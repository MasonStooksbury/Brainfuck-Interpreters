module main

fn main() {

	mut things := [1,2,3,4,5]

	println(things.last())

}